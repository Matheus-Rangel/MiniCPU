library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity registers is
    generic (
        DATA_WIDTH : integer := 16;
        ADDR_WIDTH : integer := 3
    );
    port (
        clock  : in std_logic;
        reset 	: in std_logic;
		  wren   : in std_logic;
        addr   : in std_logic_vector(ADDR_WIDTH - 1 downto 0);
        data_i : in std_logic_vector(DATA_WIDTH - 1 downto 0);
        data_o : out std_logic_vector(DATA_WIDTH - 1 downto 0)
    );
end registers;

architecture reg_arch of registers is
    type ram_t is array (0 to 2**ADDR_WIDTH - 1) of std_logic_vector(DATA_WIDTH - 1 downto 0);
    signal ram_image : ram_t := (others => x"0000");
begin
    process (clock)
    begin
        if clock'event and clock = '1' then
            data_o <= ram_image(to_integer(unsigned(addr)));
            if wren = '1' then
                ram_image(to_integer(unsigned(addr))) <= data_i;
            end if;
				if reset = '1' then
					ram_image := (others => x"0000");
        end if;
    end process;
end reg_arch;
